module d_x( 
input clk,
input go_index_in,
input signed [15:0] T,
input signed [15:0] ST,
input signed [15:0] Q,
output reg MI,
output reg MI_DONE
//output reg [3:0] state_op,
//output reg [7:0] i_op
    );
    
    parameter N = 110; //n_SV
    //corrected bias is 3.10 with accuracy 97.9%
    reg signed [150:0] b = 151'd16878005399278547787783380528615703288217; //(2**132)*bias
    reg signed [31:0] d_i [110:1]; //dual coefficients
    reg signed [31:0] x_i_1 [110:1]; //1st elements in SVs
    reg signed [31:0] x_i_2 [110:1]; //2nd elements in SVs
    reg signed [31:0] x_i_3 [110:1]; //3rd elements is SVs
    reg signed [15:0] x [3:1]; //input vector for testing
    reg x_load = 0;
    reg HALT = 0;
    reg data_load = 0; //load d_i,all x_i,x if 0
    reg [3:0] state = 0;
    reg [7:0] i = 1;
    reg signed [31:0] temp1,temp2,temp3,temp4 = 0;
    reg signed [41:0] temp6 = 0;
    reg signed [31:0] temp6_int = 0;
    reg signed [31:0] gamma = 32'd429496;//(2**32)*gamma
    reg signed [63:0] temp5 = 0;
    reg signed [200:0] temp7,temp7_9,temp7_8,temp7_7,temp7_6,temp7_5,temp7_4,temp7_3,temp7_2,temp7_1,temp7_0,temp7b;
    reg signed [250:0] temp8,temp8b = 0;
    
    
    always@(posedge clk) begin
    //state_op <= state;
    //i_op <= i;
    if ((!HALT)&&(go_index_in)) begin
    if ((!x_load)) begin
    x[1] <= T;
    x[2] <= ST;
    x[3] <= Q;
    x_load <= 1;
    end
    if (!data_load) begin
    d_i[1] <= -32'd100;
    x_i_1[1] <= 32'd372;
    x_i_2[1] <= 32'd45;
    x_i_3[1] <= 32'd36;
    d_i[2] <= -32'd100;
    x_i_1[2] <= 32'd358;
    x_i_2[2] <= 32'd42;
    x_i_3[2] <= 32'd80;
    d_i[3] <= -32'd100;
    x_i_1[3] <= -32'd147;
    x_i_2[3] <= 32'd26;
    x_i_3[3] <= 32'd56;
    d_i[4] <= -32'd100;
    x_i_1[4] <= 32'd354;
    x_i_2[4] <= 32'd42;
    x_i_3[4] <= 32'd22;
    d_i[5] <= -32'd38;
    x_i_1[5] <= 32'd473;
    x_i_2[5] <= 32'd33;
    x_i_3[5] <= 32'd64;
    d_i[6] <= -32'd100;
    x_i_1[6] <= 32'd278;
    x_i_2[6] <= 32'd45;
    x_i_3[6] <= 32'd58;
    d_i[7] <= -32'd9;
    x_i_1[7] <= -32'd66;
    x_i_2[7] <= 32'd38;
    x_i_3[7] <= 32'd20;
    d_i[8] <= -32'd50;
    x_i_1[8] <= 32'd270;
    x_i_2[8] <= 32'd40;
    x_i_3[8] <= 32'd128;
    d_i[9] <= -32'd29;
    x_i_1[9] <= -32'd80;
    x_i_2[9] <= 32'd13;
    x_i_3[9] <= 32'd67;
    d_i[10] <= -32'd100;
    x_i_1[10] <= 32'd494;
    x_i_2[10] <= 32'd29;
    x_i_3[10] <= 32'd45;
    d_i[11] <= -32'd100;
    x_i_1[11] <= 32'd478;
    x_i_2[11] <= 32'd36;
    x_i_3[11] <= 32'd41;
    d_i[12] <= -32'd100;
    x_i_1[12] <= 32'd207;
    x_i_2[12] <= 32'd44;
    x_i_3[12] <= 32'd64;
    d_i[13] <= -32'd19;
    x_i_1[13] <= 32'd404;
    x_i_2[13] <= 32'd43;
    x_i_3[13] <= 32'd85;
    d_i[14] <= -32'd94;
    x_i_1[14] <= 32'd190;
    x_i_2[14] <= 32'd41;
    x_i_3[14] <= 32'd71;
    d_i[15] <= -32'd100;
    x_i_1[15] <= 32'd94;
    x_i_2[15] <= 32'd41;
    x_i_3[15] <= 32'd82;
    d_i[16] <= -32'd55;
    x_i_1[16] <= 32'd230;
    x_i_2[16] <= 32'd41;
    x_i_3[16] <= 32'd42;
    d_i[17] <= -32'd100;
    x_i_1[17] <= 32'd172;
    x_i_2[17] <= 32'd47;
    x_i_3[17] <= 32'd46;
    d_i[18] <= -32'd29;
    x_i_1[18] <= -32'd109;
    x_i_2[18] <= 32'd41;
    x_i_3[18] <= 32'd157;
    d_i[19] <= -32'd100;
    x_i_1[19] <= 32'd360;
    x_i_2[19] <= 32'd43;
    x_i_3[19] <= 32'd62;
    d_i[20] <= -32'd100;
    x_i_1[20] <= 32'd203;
    x_i_2[20] <= 32'd40;
    x_i_3[20] <= 32'd76;
    d_i[21] <= -32'd63;
    x_i_1[21] <= 32'd438;
    x_i_2[21] <= 32'd43;
    x_i_3[21] <= 32'd65;
    d_i[22] <= -32'd100;
    x_i_1[22] <= 32'd148;
    x_i_2[22] <= 32'd44;
    x_i_3[22] <= 32'd88;
    d_i[23] <= -32'd100;
    x_i_1[23] <= 32'd258;
    x_i_2[23] <= 32'd42;
    x_i_3[23] <= 32'd77;
    d_i[24] <= -32'd100;
    x_i_1[24] <= 32'd283;
    x_i_2[24] <= 32'd49;
    x_i_3[24] <= 32'd104;
    d_i[25] <= -32'd100;
    x_i_1[25] <= 32'd254;
    x_i_2[25] <= 32'd44;
    x_i_3[25] <= 32'd24;
    d_i[26] <= -32'd96;
    x_i_1[26] <= 32'd418;
    x_i_2[26] <= 32'd45;
    x_i_3[26] <= 32'd98;
    d_i[27] <= -32'd74;
    x_i_1[27] <= 32'd142;
    x_i_2[27] <= 32'd44;
    x_i_3[27] <= 32'd52;
    d_i[28] <= -32'd54;
    x_i_1[28] <= 32'd224;
    x_i_2[28] <= 32'd42;
    x_i_3[28] <= 32'd165;
    d_i[29] <= -32'd37;
    x_i_1[29] <= -32'd202;
    x_i_2[29] <= 32'd31;
    x_i_3[29] <= 32'd124;
    d_i[30] <= -32'd100;
    x_i_1[30] <= 32'd408;
    x_i_2[30] <= 32'd49;
    x_i_3[30] <= 32'd20;
    d_i[31] <= -32'd100;
    x_i_1[31] <= 32'd204;
    x_i_2[31] <= 32'd44;
    x_i_3[31] <= 32'd31;
    d_i[32] <= -32'd1;
    x_i_1[32] <= 32'd91;
    x_i_2[32] <= 32'd39;
    x_i_3[32] <= 32'd150;
    d_i[33] <= -32'd100;
    x_i_1[33] <= 32'd192;
    x_i_2[33] <= 32'd48;
    x_i_3[33] <= 32'd33;
    d_i[34] <= -32'd2;
    x_i_1[34] <= 32'd91;
    x_i_2[34] <= 32'd39;
    x_i_3[34] <= 32'd150;
    d_i[35] <= -32'd88;
    x_i_1[35] <= -32'd93;
    x_i_2[35] <= -32'd11;
    x_i_3[35] <= 32'd183;
    d_i[36] <= -32'd100;
    x_i_1[36] <= 32'd254;
    x_i_2[36] <= 32'd44;
    x_i_3[36] <= 32'd24;
    d_i[37] <= -32'd100;
    x_i_1[37] <= 32'd254;
    x_i_2[37] <= 32'd41;
    x_i_3[37] <= 32'd56;
    d_i[38] <= -32'd2;
    x_i_1[38] <= 32'd219;
    x_i_2[38] <= 32'd42;
    x_i_3[38] <= 32'd17;
    d_i[39] <= -32'd16;
    x_i_1[39] <= 32'd129;
    x_i_2[39] <= 32'd32;
    x_i_3[39] <= 32'd185;
    d_i[40] <= -32'd11;
    x_i_1[40] <= 32'd255;
    x_i_2[40] <= 32'd40;
    x_i_3[40] <= 32'd8;
    d_i[41] <= -32'd100;
    x_i_1[41] <= 32'd452;
    x_i_2[41] <= 32'd42;
    x_i_3[41] <= 32'd55;
    d_i[42] <= -32'd40;
    x_i_1[42] <= 32'd320;
    x_i_2[42] <= 32'd42;
    x_i_3[42] <= 32'd124;
    d_i[43] <= -32'd4;
    x_i_1[43] <= 32'd336;
    x_i_2[43] <= 32'd41;
    x_i_3[43] <= -32'd26;
    d_i[44] <= -32'd100;
    x_i_1[44] <= -32'd92;
    x_i_2[44] <= 32'd28;
    x_i_3[44] <= 32'd14;
    d_i[45] <= -32'd100;
    x_i_1[45] <= 32'd316;
    x_i_2[45] <= 32'd43;
    x_i_3[45] <= 32'd56;
    d_i[46] <= -32'd100;
    x_i_1[46] <= 32'd269;
    x_i_2[46] <= 32'd55;
    x_i_3[46] <= 32'd85;
    d_i[47] <= -32'd6;
    x_i_1[47] <= 32'd386;
    x_i_2[47] <= -32'd15;
    x_i_3[47] <= 32'd26;
    d_i[48] <= -32'd100;
    x_i_1[48] <= 32'd196;
    x_i_2[48] <= 32'd61;
    x_i_3[48] <= 32'd58;
    d_i[49] <= -32'd100;
    x_i_1[49] <= -32'd86;
    x_i_2[49] <= 32'd28;
    x_i_3[49] <= 32'd85;
    d_i[50] <= -32'd100;
    x_i_1[50] <= 32'd497;
    x_i_2[50] <= 32'd39;
    x_i_3[50] <= 32'd23;
    d_i[51] <= -32'd90;
    x_i_1[51] <= 32'd74;
    x_i_2[51] <= 32'd48;
    x_i_3[51] <= 32'd57;
    d_i[52] <= -32'd100;
    x_i_1[52] <= 32'd511;
    x_i_2[52] <= 32'd46;
    x_i_3[52] <= 32'd0;
    d_i[53] <= -32'd100;
    x_i_1[53] <= 32'd193;
    x_i_2[53] <= 32'd44;
    x_i_3[53] <= 32'd43;
    d_i[54] <= -32'd70;
    x_i_1[54] <= 32'd141;
    x_i_2[54] <= 32'd55;
    x_i_3[54] <= 32'd10;
    d_i[55] <= -32'd32;
    x_i_1[55] <= 32'd124;
    x_i_2[55] <= 32'd44;
    x_i_3[55] <= 32'd115;
    d_i[56] <= 32'd100;
    x_i_1[56] <= 32'd224;
    x_i_2[56] <= 32'd46;
    x_i_3[56] <= 32'd13;
    d_i[57] <= 32'd61;
    x_i_1[57] <= 32'd238;
    x_i_2[57] <= 32'd51;
    x_i_3[57] <= 32'd143;
    d_i[58] <= 32'd25;
    x_i_1[58] <= 32'd147;
    x_i_2[58] <= 32'd24;
    x_i_3[58] <= 32'd204;
    d_i[59] <= 32'd100;
    x_i_1[59] <= 32'd176;
    x_i_2[59] <= 32'd46;
    x_i_3[59] <= 32'd77;
    d_i[60] <= 32'd78;
    x_i_1[60] <= 32'd446;
    x_i_2[60] <= 32'd51;
    x_i_3[60] <= 32'd49;
    d_i[61] <= 32'd100;
    x_i_1[61] <= -32'd92;
    x_i_2[61] <= 32'd31;
    x_i_3[61] <= 32'd17;
    d_i[62] <= 32'd29;
    x_i_1[62] <= 32'd238;
    x_i_2[62] <= -32'd27;
    x_i_3[62] <= 32'd69;
    d_i[63] <= 32'd100;
    x_i_1[63] <= 32'd170;
    x_i_2[63] <= 32'd50;
    x_i_3[63] <= 32'd53;
    d_i[64] <= 32'd68;
    x_i_1[64] <= 32'd471;
    x_i_2[64] <= 32'd49;
    x_i_3[64] <= 32'd48;
    d_i[65] <= 32'd12;
    x_i_1[65] <= -32'd148;
    x_i_2[65] <= 32'd44;
    x_i_3[65] <= 32'd97;
    d_i[66] <= 32'd100;
    x_i_1[66] <= 32'd233;
    x_i_2[66] <= 32'd45;
    x_i_3[66] <= 32'd53;
    d_i[67] <= 32'd100;
    x_i_1[67] <= 32'd356;
    x_i_2[67] <= 32'd47;
    x_i_3[67] <= 32'd72;
    d_i[68] <= 32'd100;
    x_i_1[68] <= 32'd165;
    x_i_2[68] <= 32'd47;
    x_i_3[68] <= 32'd45;
    d_i[69] <= 32'd21;
    x_i_1[69] <= 32'd49;
    x_i_2[69] <= 32'd51;
    x_i_3[69] <= 32'd95;
    d_i[70] <= 32'd100;
    x_i_1[70] <= 32'd138;
    x_i_2[70] <= 32'd47;
    x_i_3[70] <= 32'd70;
    d_i[71] <= 32'd89;
    x_i_1[71] <= 32'd279;
    x_i_2[71] <= 32'd51;
    x_i_3[71] <= 32'd83;
    d_i[72] <= 32'd4;
    x_i_1[72] <= 32'd255;
    x_i_2[72] <= 32'd49;
    x_i_3[72] <= 32'd34;
    d_i[73] <= 32'd2;
    x_i_1[73] <= 32'd185;
    x_i_2[73] <= 32'd42;
    x_i_3[73] <= 32'd215;
    d_i[74] <= 32'd100;
    x_i_1[74] <= -32'd86;
    x_i_2[74] <= 32'd28;
    x_i_3[74] <= 32'd85;
    d_i[75] <= 32'd1;
    x_i_1[75] <= -32'd252;
    x_i_2[75] <= 32'd37;
    x_i_3[75] <= 32'd95;
    d_i[76] <= 32'd100;
    x_i_1[76] <= 32'd258;
    x_i_2[76] <= 32'd48;
    x_i_3[76] <= 32'd33;
    d_i[77] <= 32'd69;
    x_i_1[77] <= 32'd238;
    x_i_2[77] <= 32'd43;
    x_i_3[77] <= 32'd115;
    d_i[78] <= 32'd7;
    x_i_1[78] <= -32'd159;
    x_i_2[78] <= 32'd24;
    x_i_3[78] <= 32'd135;
    d_i[79] <= 32'd100;
    x_i_1[79] <= 32'd404;
    x_i_2[79] <= 32'd48;
    x_i_3[79] <= 32'd50;
    d_i[80] <= 32'd20;
    x_i_1[80] <= 32'd338;
    x_i_2[80] <= 32'd49;
    x_i_3[80] <= 32'd60;
    d_i[81] <= 32'd100;
    x_i_1[81] <= 32'd367;
    x_i_2[81] <= 32'd46;
    x_i_3[81] <= 32'd25;
    d_i[82] <= 32'd100;
    x_i_1[82] <= 32'd284;
    x_i_2[82] <= 32'd46;
    x_i_3[82] <= 32'd66;
    d_i[83] <= 32'd100;
    x_i_1[83] <= 32'd210;
    x_i_2[83] <= 32'd47;
    x_i_3[83] <= 32'd47;
    d_i[84] <= 32'd40;
    x_i_1[84] <= 32'd391;
    x_i_2[84] <= -32'd24;
    x_i_3[84] <= 32'd50;
    d_i[85] <= 32'd47;
    x_i_1[85] <= -32'd194;
    x_i_2[85] <= 32'd19;
    x_i_3[85] <= 32'd83;
    d_i[86] <= 32'd100;
    x_i_1[86] <= 32'd389;
    x_i_2[86] <= 32'd47;
    x_i_3[86] <= 32'd94;
    d_i[87] <= 32'd100;
    x_i_1[87] <= 32'd91;
    x_i_2[87] <= 32'd48;
    x_i_3[87] <= 32'd49;
    d_i[88] <= 32'd100;
    x_i_1[88] <= 32'd186;
    x_i_2[88] <= 32'd49;
    x_i_3[88] <= 32'd26;
    d_i[89] <= 32'd100;
    x_i_1[89] <= 32'd440;
    x_i_2[89] <= 32'd46;
    x_i_3[89] <= 32'd44;
    d_i[90] <= 32'd100;
    x_i_1[90] <= 32'd501;
    x_i_2[90] <= 32'd40;
    x_i_3[90] <= 32'd25;
    d_i[91] <= 32'd82;
    x_i_1[91] <= 32'd348;
    x_i_2[91] <= 32'd47;
    x_i_3[91] <= 32'd26;
    d_i[92] <= 32'd100;
    x_i_1[92] <= 32'd177;
    x_i_2[92] <= 32'd53;
    x_i_3[92] <= 32'd29;
    d_i[93] <= 32'd100;
    x_i_1[93] <= 32'd202;
    x_i_2[93] <= 32'd45;
    x_i_3[93] <= 32'd80;
    d_i[94] <= 32'd82;
    x_i_1[94] <= 32'd94;
    x_i_2[94] <= 32'd46;
    x_i_3[94] <= 32'd90;
    d_i[95] <= 32'd100;
    x_i_1[95] <= 32'd238;
    x_i_2[95] <= 32'd45;
    x_i_3[95] <= 32'd71;
    d_i[96] <= 32'd100;
    x_i_1[96] <= 32'd509;
    x_i_2[96] <= 32'd32;
    x_i_3[96] <= 32'd14;
    d_i[97] <= 32'd18;
    x_i_1[97] <= -32'd54;
    x_i_2[97] <= -32'd52;
    x_i_3[97] <= 32'd167;
    d_i[98] <= 32'd76;
    x_i_1[98] <= 32'd507;
    x_i_2[98] <= 32'd29;
    x_i_3[98] <= 32'd28;
    d_i[99] <= 32'd73;
    x_i_1[99] <= -32'd107;
    x_i_2[99] <= -32'd6;
    x_i_3[99] <= 32'd197;
    d_i[100] <= 32'd100;
    x_i_1[100] <= 32'd272;
    x_i_2[100] <= 32'd43;
    x_i_3[100] <= 32'd79;
    d_i[101] <= 32'd94;
    x_i_1[101] <= 32'd255;
    x_i_2[101] <= 32'd49;
    x_i_3[101] <= 32'd34;
    d_i[102] <= 32'd100;
    x_i_1[102] <= 32'd330;
    x_i_2[102] <= 32'd46;
    x_i_3[102] <= 32'd38;
    d_i[103] <= 32'd55;
    x_i_1[103] <= -32'd111;
    x_i_2[103] <= 32'd28;
    x_i_3[103] <= 32'd115;
    d_i[104] <= 32'd100;
    x_i_1[104] <= 32'd319;
    x_i_2[104] <= 32'd48;
    x_i_3[104] <= 32'd120;
    d_i[105] <= 32'd42;
    x_i_1[105] <= 32'd118;
    x_i_2[105] <= 32'd48;
    x_i_3[105] <= 32'd95;
    d_i[106] <= 32'd100;
    x_i_1[106] <= 32'd471;
    x_i_2[106] <= 32'd31;
    x_i_3[106] <= 32'd87;
    d_i[107] <= 32'd39;
    x_i_1[107] <= 32'd457;
    x_i_2[107] <= 32'd56;
    x_i_3[107] <= 32'd6;
    d_i[108] <= 32'd72;
    x_i_1[108] <= -32'd120;
    x_i_2[108] <= 32'd21;
    x_i_3[108] <= 32'd34;
    d_i[109] <= 32'd5;
    x_i_1[109] <= 32'd250;
    x_i_2[109] <= -32'd35;
    x_i_3[109] <= 32'd41;
    d_i[110] <= 32'd100;
    x_i_1[110] <= 32'd219;
    x_i_2[110] <= 32'd45;
    x_i_3[110] <= 32'd58;
    data_load <= 1;
    end
    else begin
    if (i <= 110) begin
        if (state == 5) begin
            i <= i + 1;
            temp8b <= temp8b + temp8;//this is origional sigma di*K(x,xi)*(2**132)
            state <= 1;
        end
        else state <= state + 1;
    end
    else begin
        MI <= ((temp8b + b)>=0)?1:0;
        MI_DONE <= 1;
        HALT <= 1;
        i <= 110;
        state <= 0;
    end
    end
    end
    end
    
    
    always@(*) begin
    if ((!HALT)&&(i >= 1)&&(i <= 110)&&(data_load == 1)&&(state > 0)&&(go_index_in)) begin
        case(state)
        1: begin
           temp1 = (x[1] - x_i_1[i])*(x[1] - x_i_1[i]);
           temp2 = (x[2] - x_i_2[i])*(x[2] - x_i_2[i]);
           temp3 = (x[3] - x_i_3[i])*(x[3] - x_i_3[i]);
           temp4 = temp1 + temp2 + temp3;
           temp5 = 0;
           temp6 = 0;
           temp6_int = 0;
           temp7 = 0;
           temp7_0 = 0;
           temp7_1 = 0;
           temp7_2 = 0;
           temp7_3 = 0;
           temp7_4 = 0;
           temp7_5 = 0;
           temp7_6 = 0;
           temp7_7 = 0;
           temp7_8 = 0;
           temp7_9 = 0;
           temp7b = 0;
           temp8 = 0;
           end
        2: begin
           temp1 = (x[1] - x_i_1[i])*(x[1] - x_i_1[i]);
           temp2 = (x[2] - x_i_2[i])*(x[2] - x_i_2[i]);
           temp3 = (x[3] - x_i_3[i])*(x[3] - x_i_3[i]);
           temp4 = temp1 + temp2 + temp3;
           temp5 = temp4*gamma;
           temp6 = temp5[63:22];
           temp6_int = temp5[63:32];
           temp7 = 0;
           temp7_0 = 0;
           temp7_1 = 0;
           temp7_2 = 0;
           temp7_3 = 0;
           temp7_4 = 0;
           temp7_5 = 0;
           temp7_6 = 0;
           temp7_7 = 0;
           temp7_8 = 0;
           temp7_9 = 0;
           temp7b = 0;
           temp8 = 0;
           end
        3: begin
           temp1 = (x[1] - x_i_1[i])*(x[1] - x_i_1[i]);
           temp2 = (x[2] - x_i_2[i])*(x[2] - x_i_2[i]);
           temp3 = (x[3] - x_i_3[i])*(x[3] - x_i_3[i]);
           temp4 = temp1 + temp2 + temp3;
           temp5 = temp4*gamma;
           temp6 = temp5[63:22];
           temp6_int = temp5[63:32];
           if (temp6_int < 11) begin
           temp7 = (temp6_int==0)?64'd4294967296:0;
           temp7 = (temp6_int==1)?64'd1580030168:0;
           temp7 = (temp6_int==2)?64'd581260615:0;
           temp7 = (temp6_int==3)?64'd213833830:0;
           temp7 = (temp6_int==4)?64'd78665070:0;
           temp7 = (temp6_int==5)?64'd28939262:0;
           temp7 = (temp6_int==6)?64'd10646159:0;
           temp7 = (temp6_int==7)?64'd3916503:0;
           temp7 = (temp6_int==8)?64'd1440801:0;
           temp7 = (temp6_int==9)?64'd530041:0;
           temp7 = (temp6_int==10)?64'd194991:0;
           end
           else temp7 = 0;
           
           temp7_9 = temp6[9]?(temp7*621):(temp7<<10);
           temp7_8 = temp6[8]?(temp7_9*797):(temp7_9<<10);
           temp7_7 = temp6[7]?(temp7_8*904):(temp7_8<<10);
           temp7_6 = temp6[6]?(temp7_7*962):(temp7_7<<10);
           temp7_5 = temp6[5]?(temp7_6*992):(temp7_6<<10);
           temp7_4 = temp6[4]?(temp7_5*1008):(temp7_5<<10);
           temp7_3 = temp6[3]?(temp7_4*1016):(temp7_4<<10);
           temp7_2 = temp6[2]?(temp7_3*1020):(temp7_3<<10);
           temp7_1 = temp6[1]?(temp7_2*1022):(temp7_2<<10);
           temp7_0 = temp6[0]?(temp7_1*1023):(temp7_1<<10);
           
           temp7b = 0;
           temp8 = 0;
           end
        4: begin
           temp1 = (x[1] - x_i_1[i])*(x[1] - x_i_1[i]);
           temp2 = (x[2] - x_i_2[i])*(x[2] - x_i_2[i]);
           temp3 = (x[3] - x_i_3[i])*(x[3] - x_i_3[i]);
           temp4 = temp1 + temp2 + temp3;
           temp5 = temp4*gamma;
           temp6 = temp5[63:22];
           temp6_int = temp5[63:32];
           if (temp6_int < 11) begin
           temp7 = (temp6_int==0)?64'd4294967296:0;
           temp7 = (temp6_int==1)?64'd1580030168:0;
           temp7 = (temp6_int==2)?64'd581260615:0;
           temp7 = (temp6_int==3)?64'd213833830:0;
           temp7 = (temp6_int==4)?64'd78665070:0;
           temp7 = (temp6_int==5)?64'd28939262:0;
           temp7 = (temp6_int==6)?64'd10646159:0;
           temp7 = (temp6_int==7)?64'd3916503:0;
           temp7 = (temp6_int==8)?64'd1440801:0;
           temp7 = (temp6_int==9)?64'd530041:0;
           temp7 = (temp6_int==10)?64'd194991:0;
           end
           else temp7 = 0;
           
           temp7_9 = temp6[9]?(temp7*621):(temp7<<10);
           temp7_8 = temp6[8]?(temp7_9*797):(temp7_9<<10);
           temp7_7 = temp6[7]?(temp7_8*904):(temp7_8<<10);
           temp7_6 = temp6[6]?(temp7_7*962):(temp7_7<<10);
           temp7_5 = temp6[5]?(temp7_6*992):(temp7_6<<10);
           temp7_4 = temp6[4]?(temp7_5*1008):(temp7_5<<10);
           temp7_3 = temp6[3]?(temp7_4*1016):(temp7_4<<10);
           temp7_2 = temp6[2]?(temp7_3*1020):(temp7_3<<10);
           temp7_1 = temp6[1]?(temp7_2*1022):(temp7_2<<10);
           temp7_0 = temp6[0]?(temp7_1*1023):(temp7_1<<10);
           temp7b = temp7_0*d_i[i];
           temp8 = 0;
           end
        5: begin
           temp1 = (x[1] - x_i_1[i])*(x[1] - x_i_1[i]);
           temp2 = (x[2] - x_i_2[i])*(x[2] - x_i_2[i]);
           temp3 = (x[3] - x_i_3[i])*(x[3] - x_i_3[i]);
           temp4 = temp1 + temp2 + temp3;
           temp5 = temp4*gamma;
           temp6 = temp5[63:22];
           temp6_int = temp5[63:32];
           if (temp6_int < 11) begin
           temp7 = (temp6_int==0)?64'd4294967296:0;
           temp7 = (temp6_int==1)?64'd1580030168:0;
           temp7 = (temp6_int==2)?64'd581260615:0;
           temp7 = (temp6_int==3)?64'd213833830:0;
           temp7 = (temp6_int==4)?64'd78665070:0;
           temp7 = (temp6_int==5)?64'd28939262:0;
           temp7 = (temp6_int==6)?64'd10646159:0;
           temp7 = (temp6_int==7)?64'd3916503:0;
           temp7 = (temp6_int==8)?64'd1440801:0;
           temp7 = (temp6_int==9)?64'd530041:0;
           temp7 = (temp6_int==10)?64'd194991:0;
           end
           else temp7 = 0;
           
           temp7_9 = temp6[9]?(temp7*621):(temp7<<10);
           temp7_8 = temp6[8]?(temp7_9*797):(temp7_9<<10);
           temp7_7 = temp6[7]?(temp7_8*904):(temp7_8<<10);
           temp7_6 = temp6[6]?(temp7_7*962):(temp7_7<<10);
           temp7_5 = temp6[5]?(temp7_6*992):(temp7_6<<10);
           temp7_4 = temp6[4]?(temp7_5*1008):(temp7_5<<10);
           temp7_3 = temp6[3]?(temp7_4*1016):(temp7_4<<10);
           temp7_2 = temp6[2]?(temp7_3*1020):(temp7_3<<10);
           temp7_1 = temp6[1]?(temp7_2*1022):(temp7_2<<10);
           temp7_0 = temp6[0]?(temp7_1*1023):(temp7_1<<10);
           temp7b = temp7_0*d_i[i];
           temp8 = temp7b;
           end
        default: begin
                 temp1 = 0;
                 temp2 = 0;
                 temp3 = 0;
                 temp4 = 0;
                 temp5 = 0;
                 temp6 = 0;
                 temp6_int = 0;
                 temp7 = 0;
                 temp7_0 = 0;
                 temp7_1 = 0;
                 temp7_2 = 0;
                 temp7_3 = 0;
                 temp7_4 = 0;
                 temp7_5 = 0;
                 temp7_6 = 0;
                 temp7_7 = 0;
                 temp7_8 = 0;
                 temp7_9 = 0;
                 temp7b = 0;
                 temp8 = 0;
                 end
        endcase
    end
    end
    
endmodule
